/home/cc/eecs151/fa23/class/eecs151-aeq/asic_labs_fa23/lab6/build/tech-sky130-cache/sky130_ef_io.lef